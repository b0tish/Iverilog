module xorgate(a,b,out);

input a,b;
output out;
xor a1(out,a,b);

endmodule
