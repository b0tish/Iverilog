module orgate(a,b,out);

input a,b;
output out;
or a1(out,a,b);

endmodule
