module andgate(a,b,out);

input a,b;
output out;
and a1(out,a,b);

endmodule
