module nandgate(a,b,out);

input a,b;
output out;
nand a1(out,a,b);

endmodule
